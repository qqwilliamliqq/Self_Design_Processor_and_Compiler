module inst_rom #(parameter A=12, W=9) (
  input		   [A-1:0] InstAddress,
  output logic [W-1:0] InstOut
  );
  
  logic [W-1:0] inst_rom[2**(A)];
  always_comb begin
    InstOut = inst_rom[InstAddress];
  end

  initial begin
	$readmemb("machine_code.txt", inst_rom);
	//$display("%s", inst_rom[0]);
  end

endmodule